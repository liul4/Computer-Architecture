library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Memory32Bit is
Port (address : in std_logic_vector(31 downto 0);
write_data : in std_logic_vector(31 downto 0);
write_enable : in std_logic;
clock : in std_logic;
read_data : out std_logic_vector(31 downto 0));
end Memory32Bit;

architecture Behavioral of Memory32Bit is
type mem_array is array(0 to 511) of std_logic_vector(31 downto 0); 
signal data_mem : mem_array := (
X"00000000", X"00000001", X"00000002",X"00000003", X"00000004", X"00000005", X"00000006",X"00000007",
X"00000008", X"00000009", 
X"0000000A",X"0000000B", X"0000000C", X"0000000D", X"0000000E",X"0000000F",
X"00000010", X"00000011", X"00000012",X"00000013", X"00000014", X"00000015", X"00000016",X"00000017",
X"00000018", X"00000019", X"0000001A",X"0000001B", X"0000001C", X"0000001D", X"0000001E",X"0000001F",
X"00000020", X"00000021", X"00000022",X"00000023", X"00000024", X"00000005", X"00000026",X"00000027",
X"00000028", X"00000029", X"0000002A",X"0000002B", X"0000002C", X"0000002D", X"0000002E",X"0000002F",
X"00000030", X"00000031", X"00000032",X"00000033",
X"00000034", X"00000035", X"00000036",X"00000037",
X"00000038", X"00000039", X"0000003A",X"0000003B", X"0000003C", X"0000003D", X"0000003E",X"0000003F",
X"00000040", X"00000041", X"00000042",X"00000043", X"00000044", X"00000045", X"00000046",X"00000047",
X"00000048", X"00000049", X"0000004A",X"0000004B", X"0000004C", X"0000004D", X"0000004E",X"0000004F",
X"00000050", X"00000051", X"00000052",X"00000053", X"00000054", X"00000055", X"00000056",X"00000057",
X"00000058", X"00000059", X"0000005A",X"0000005B", X"0000005C", X"0000005D", X"0000005E",X"0000005F",
X"00000060", X"00000061", X"00000062",X"00000063", X"00000064", X"00000065", X"00000066",X"00000067",
X"00000068", X"00000069", X"0000006A",X"0000006B", X"0000006C", X"0000006D", X"0000006E",X"0000006F",
X"00000070", X"00000071", X"00000072",X"00000073", X"00000074", X"00000075", X"00000076",X"00000077",
X"00000078", X"00000079", X"0000007A",X"0000007B", X"0000007C", X"0000007D", X"0000007E",X"0000007F",
X"00000080", X"00000081", X"00000082",X"00000083", X"00000084", X"00000085", X"00000086",X"00000087",
X"00000088", X"00000089", X"0000008A",X"0000008B", X"0000008C", X"0000008D", X"0000008E",X"0000008F",
X"00000090", X"00000091", X"00000092",X"00000093", X"00000094", X"00000095", X"00000096",X"00000097",
X"00000098", X"00000099", X"0000009A",X"0000009B", X"0000009C", X"0000009D", X"0000009E",X"0000009F",
X"000000A0", X"000000A1", X"000000A2",X"000000A3", X"000000A4", X"000000A5", X"000000A6",X"000000A7",
X"000000A8", X"000000A9", X"000000AA",X"000000AB", X"000000AC", X"000000AD", X"000000AE",X"000000AF",
X"000000B0", X"000000B1", X"000000B2",X"000000B3", X"000000B4", X"000000B5", X"000000B6",X"000000B7",
X"000000B8", X"000000B9", X"000000BA",X"000000BB", X"000000BC", X"000000BD", X"000000BE",X"000000BF",
X"000000C0", X"000000C1", X"000000C2",X"000000C3", X"000000C4", X"000000C5", X"000000C6",X"000000C7",
X"000000C8", X"000000C9", X"000000CA",X"000000CB", X"000000CC", X"000000CD", X"000000CE",X"000000CF",
X"000000D0", X"000000D1", X"000000D2",X"000000D3", X"000000D4", X"000000D5", X"000000D6",X"000000D7",
X"000000D8", X"000000D9", X"000000DA",X"000000DB", X"000000DC", X"000000DD", X"000000DE",X"000000DF",
X"000000E0", X"000000E1", X"000000E2",X"000000E3", X"000000E4", X"000000E5", X"000000E6",X"000000E7",
X"000000E8", X"000000E9", X"000000EA",X"000000EB", X"000000EC", X"000000ED", X"000000EE",X"000000EF",
X"000000F0", X"000000F1", X"000000F2",X"000000F3", X"000000F4", X"000000F5", X"000000F6",X"000000F7",
X"000000F8", X"000000F9", X"000000FA",X"000000FB", X"000000FC", X"000000FD", X"000000FE",X"000000FF",
X"00000100", X"00000101", X"00000102",X"00000103", X"00000104", X"00000105", X"00000106",X"00000107",
X"00000108", X"00000109", X"0000010A",X"0000010B", X"0000010C", X"0000010D", X"0000010E",X"0000010F",
X"00000110", X"00000111", X"00000112",X"00000113", X"00000114", X"00000115", X"00000116",X"00000117",
X"00000118", X"00000119", X"0000011A",X"0000011B", X"0000011C", X"0000011D", X"0000011E",X"0000011F",
X"00000120", X"00000121", X"00000122",X"00000123", X"00000124", X"00000105", X"00000126",X"00000127",
X"00000128", X"00000129", X"0000012A",X"0000012B", X"0000012C", X"0000012D", X"0000012E",X"0000012F",
X"00000130", X"00000131", X"00000132",X"00000133", X"00000134", X"00000135", X"00000136",X"00000137",
X"00000138", X"00000139", X"0000013A",X"0000013B", X"0000013C", X"0000013D", X"0000013E",X"0000013F",
X"00000140", X"00000141", X"00000142",X"00000143", X"00000144", X"00000145", X"00000146",X"00000147",
X"00000148", X"00000149", X"0000014A",X"0000014B", X"0000014C", X"0000014D", X"0000014E",X"0000014F",
X"00000150", X"00000151", X"00000152",X"00000153", X"00000154", X"00000155", X"00000156",X"00000157",
X"00000158", X"00000159", X"0000015A",X"0000015B", X"0000015C", X"0000015D", X"0000015E",X"0000015F",
X"00000160", X"00000161", X"00000162",X"00000163", X"00000164", X"00000165", X"00000166",X"00000167",
X"00000168", X"00000169", X"0000016A",X"0000016B", X"0000016C", X"0000016D", X"0000016E",X"0000016F",
X"00000170", X"00000171", X"00000172",X"00000173", X"00000174", X"00000175", X"00000176",X"00000177",
X"00000178", X"00000179", X"0000017A",X"0000017B", X"0000017C", X"0000017D", X"0000017E",X"0000017F",
X"00000180", X"00000181", X"00000182",X"00000183", X"00000184", X"00000185", X"00000186",X"00000187",
X"00000188", X"00000189", X"0000018A",X"0000018B", X"0000018C", X"0000018D", X"0000018E",X"0000018F",
X"00000190", X"00000191", X"00000192",X"00000193", X"00000194", X"00000195", X"00000196",X"00000197",
X"00000198", X"00000199", X"0000019A",X"0000019B", X"0000019C", X"0000019D", X"0000019E",X"0000019F",
X"000001A0", X"000001A1", X"000001A2",X"000001A3", X"000001A4", X"000001A5", X"000001A6",X"000001A7",
X"000001A8", X"000001A9", X"000001AA",X"000001AB", X"000001AC", X"000001AD", X"000001AE",X"000001AF",
X"000001B0", X"000001B1", X"000001B2",X"000001B3", X"000001B4", X"000001B5", X"000001B6",X"000001B7",
X"000001B8", X"000001B9", X"000001BA",X"000001BB", X"000001BC", X"000001BD", X"000001BE",X"000001BF",
X"000001C0", X"000001C1", X"000001C2",X"000001C3", X"000001C4", X"000001C5", X"000001C6",X"000001C7",
X"000001C8", X"000001C9", X"000001CA",X"000001CB", X"000001CC", X"000001CD", X"000001CE",X"000001CF",
X"000001D0", X"000001D1", X"000001D2",X"000001D3", X"000001D4", X"000001D5", X"000001D6",X"000001D7",
X"000001D8", X"000001D9", X"000001DA",X"000001DB", X"000001DC", X"000001DD", X"000001DE",X"000001DF",
X"000001E0", X"000001E1", X"000001E2",X"000001E3", X"000001E4", X"000001E5", X"000001E6",X"000001E7",
X"000001E8", X"000001E9", X"000001EA",X"000001EB", X"000001EC", X"000001ED", X"000001EE",X"000001EF",
X"000001F0", X"000001F1", X"000001F2",X"000001F3", X"000001F4", X"000001F5", X"000001F6",X"000001F7",
X"000001F8", X"000001F9", X"000001FA",X"000001FB", X"000001FC", X"000001FD", X"000001FE",X"000001FF"
); 
begin
mem_process: process(clock)
begin
if(rising_edge(clock)) then
if(write_enable='1') then
data_mem(to_integer(unsigned(address))) <= write_data after 2ns;
end if;
end if;
end process;
read_data <= data_mem(to_integer(unsigned(address))) after 2ns;
end Behavioral;
