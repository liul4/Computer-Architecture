library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
entity Memory32Bit_tb is
--  Port ( );
end Memory32Bit_tb;

architecture Behavioral of Memory32Bit_tb is
COMPONENT Memory32Bit
Port (address : in std_logic_vector(31 downto 0);
write_data : in std_logic_vector(31 downto 0);
write_enable : in std_logic;
clock : in std_logic;
read_data : out std_logic_vector(31 downto 0));
END COMPONENT;
--Inputs
signal address : std_logic_vector(31 downto 0) := (others => '0');
signal write_data : std_logic_vector(31 downto 0) := (others => '0');
signal write_enable : std_logic := '0';
signal clock : std_logic := '0';
--Outputs
signal read_data : std_logic_vector(31 downto 0);
--constant
constant PERIOD : time := 20ns;
begin
uut: Memory32Bit PORT MAP (
  address=>address,
  write_data=>write_data,
  write_enable=>write_enable,
  clock=>clock,
  read_data=>read_data
);
clock <= not clock after PERIOD/2;
stim_proc: process
  begin
  write_enable<='0';
  address<=X"00000000";
  write_data<=X"00000052"; 
  wait until clock'event and clock='1';
  address<=X"00000001";
  write_data<=X"00000053";
  wait until clock'event and clock='1';
  address<=X"00000002";
  write_data<= X"00000054";
  wait until clock'event and clock='1';
  address<=X"00000003";
  write_data<=X"00000055";
  wait until clock'event and clock='1';
  address<=X"00000004";
  write_data<= X"00000056";
  wait until clock'event and clock='1';
  address<=X"00000005";
  write_data<= X"00000057";
  wait until clock'event and clock='1';
  address<=X"00000006";
  write_data<= X"00000058";
  wait until clock'event and clock='1';
  address<=X"00000007";
  write_data<=X"00000059";
  wait until clock'event and clock='1';
  address<=X"00000008";
  write_data<=X"00000060";
  wait until clock'event and clock='1';
  address<=X"00000009";
  write_data<= X"00000061";
  wait until clock'event and clock='1';
  address<=X"0000000A";
  write_data<= X"00000062";
  wait until clock'event and clock='1';
  address<=X"0000000B";
  write_data<=X"00000063";
  wait until clock'event and clock='1';
  address<=X"0000000C";
  write_data<= X"00000064";
  wait until clock'event and clock='1';
  address<=X"0000000D";
  write_data<= X"00000065";
  wait until clock'event and clock='1';
  address<=X"0000000E";
  write_data<= X"00000066";
  wait until clock'event and clock='1';
  address<=X"0000000F";
  write_data<=X"00000067";
  wait until clock'event and clock='1';
  address<=X"00000010";
  write_data<= X"00000068";
  wait until clock'event and clock='1';
  address<=X"00000011";
  write_data<= X"00000069";
  wait until clock'event and clock='1';
  address<=X"00000012";
  write_data<=X"00000070";
  wait until clock'event and clock='1';
  address<=X"00000013";
  write_data<= X"00000071";
  wait until clock'event and clock='1';
  address<=X"00000014";
  write_data<= X"00000072";
  wait until clock'event and clock='1';
  address<=X"00000015";
  write_data<= X"00000073";
  wait until clock'event and clock='1';
  address<=X"00000016";
  write_data<=X"00000074";
  wait until clock'event and clock='1';
  address<=X"00000017";
  write_data<= X"00000065";
  wait until clock'event and clock='1';
  address<=X"00000018";
  write_data<= X"00000066";
  wait until clock'event and clock='1';
  address<=X"00000019";
  write_data<=X"00000067";
  wait until clock'event and clock='1';
  address<=X"0000001A";
  write_data<= X"00000068";
  wait until clock'event and clock='1';
  address<=X"0000001B";
  write_data<= X"00000069";
  wait until clock'event and clock='1';
  address<=X"0000001C";
  write_data<=X"00000080";
  wait until clock'event and clock='1';
  address<=X"0000001D";
  write_data<= X"00000081";
  wait until clock'event and clock='1';
  address<=X"0000001E";
  write_data<= X"00000082";
  wait until clock'event and clock='1';
  address<=X"0000001F";
  write_data<= X"00000083";
  wait until clock'event and clock='1';
  address<=X"00000020";
  write_data<=X"00000084";
  wait until clock'event and clock='1';
  address<=X"00000021";
  write_data<= X"00000085";
  wait until clock'event and clock='1';
  address<=X"00000022";
  write_data<= X"00000086";
  wait until clock'event and clock='1';
  address<=X"00000023";
  write_data<=X"00000087";
  wait until clock'event and clock='1';
  address<=X"00000024";
  write_data<= X"00000088";
  wait until clock'event and clock='1';
  address<=X"00000025";
  write_data<= X"00000089";
  wait until clock'event and clock='1';
  address<=X"00000026";
  write_data<=X"00000090";
  wait until clock'event and clock='1';
  address<=X"00000027";
  write_data<= X"00000091";
  wait until clock'event and clock='1';
  address<=X"00000028";
  write_data<= X"00000092";
  wait until clock'event and clock='1';
  address<=X"00000029";
  write_data<= X"00000093";
  wait until clock'event and clock='1';
  address<=X"0000002A";
  write_data<=X"00000094";
  wait until clock'event and clock='1';
  address<=X"0000002B";
  write_data<= X"00000095";
  wait until clock'event and clock='1';
  address<=X"0000002C";
  write_data<= X"00000096";
  wait until clock'event and clock='1';
  address<=X"0000002D";
  write_data<=X"00000097";
  wait until clock'event and clock='1';
  address<=X"0000002E";
  write_data<= X"00000098";
  wait until clock'event and clock='1';
  address<=X"0000002F";
  write_data<= X"00000099";
  wait until clock'event and clock='1';
  address<=X"00000030";
  write_data<=X"00000100";
  wait until clock'event and clock='1';
  address<=X"00000031";
  write_data<= X"00000101";
  wait until clock'event and clock='1';
  address<=X"00000032";
  write_data<= X"00000102";
  wait until clock'event and clock='1';
  address<=X"00000033";
  write_data<= X"00000103";
  wait until clock'event and clock='1';
  address<=X"00000034";
  write_data<=X"00000104";
  wait until clock'event and clock='1';
  address<=X"00000035";
  write_data<= X"00000105";
  wait until clock'event and clock='1';
  address<=X"00000036";
  write_data<= X"00000106";
  wait until clock'event and clock='1';
  address<=X"00000037";
  write_data<=X"00000107";
  wait until clock'event and clock='1';
  address<=X"00000038";
  write_data<= X"00000108";
  wait until clock'event and clock='1';
  address<=X"00000039";
  write_data<= X"00000109";
  wait until clock'event and clock='1';
  address<=X"0000003A";
  write_data<=X"00000110";
  wait until clock'event and clock='1';
  address<=X"0000003B";
  write_data<= X"00000111";
  wait until clock'event and clock='1';
  address<=X"0000003C";
  write_data<= X"00000112";
  wait until clock'event and clock='1';
  address<=X"0000003D";
  write_data<= X"00000113";
  wait until clock'event and clock='1';
  address<=X"0000003E";
  write_data<=X"00000114";
  wait until clock'event and clock='1';
  address<=X"0000003F";
  write_data<= X"00000115";
  wait until clock'event and clock='1';
  address<=X"00000040";
  write_data<= X"00000116";
  wait until clock'event and clock='1';
  address<=X"00000041";
  write_data<=X"00000117";
  wait until clock'event and clock='1';
  address<=X"00000042";
  write_data<= X"00000118";
  wait until clock'event and clock='1';
  address<=X"00000043";
  write_data<= X"00000119";
  wait until clock'event and clock='1';
  address<=X"00000044";
  write_data<=X"00000120";
  wait until clock'event and clock='1';
  address<=X"00000045";
  write_data<= X"00000121";
  wait until clock'event and clock='1';
  address<=X"00000046";
  write_data<= X"00000122";
  wait until clock'event and clock='1';
  address<=X"00000047";
  write_data<= X"00000123";
  wait until clock'event and clock='1';
  address<=X"00000048";
  write_data<=X"00000124";
  wait until clock'event and clock='1';
  address<=X"00000049";
  write_data<= X"00000125";
  wait until clock'event and clock='1';
  address<=X"0000004A";
  write_data<= X"00000126";
  wait until clock'event and clock='1';
  address<=X"0000004B";
  write_data<=X"00000127";
  wait until clock'event and clock='1';
  address<=X"0000004C";
  write_data<= X"00000128";
  wait until clock'event and clock='1';
  address<=X"0000004D";
  write_data<= X"00000129";
  wait until clock'event and clock='1';
  address<=X"0000004E";
  write_data<=X"00000130";
  wait until clock'event and clock='1';
  address<=X"0000004F";
  write_data<= X"00000131";
  wait until clock'event and clock='1';
  address<=X"00000050";
  write_data<= X"00000132";
  wait until clock'event and clock='1';
  address<=X"00000051";
  write_data<= X"00000133";
  wait until clock'event and clock='1';
  address<=X"00000052";
  write_data<=X"00000134";
  wait until clock'event and clock='1';
  address<=X"00000053";
  write_data<=X"00000135";
  wait until clock'event and clock='1';
  address<=X"00000054";
  write_data<= X"00000136";
  wait until clock'event and clock='1';
  address<=X"00000055";
  write_data<=X"00000137";
  wait until clock'event and clock='1';
  address<=X"00000056";
  write_data<= X"00000138";
  wait until clock'event and clock='1';
  address<=X"00000057";
  write_data<= X"00000139";
  wait until clock'event and clock='1';
  address<=X"00000058";
  write_data<=X"00000140";
  wait until clock'event and clock='1';
  address<=X"00000059";
  write_data<= X"00000141";
  wait until clock'event and clock='1';
  address<=X"0000005A";
  write_data<= X"00000142";
  wait until clock'event and clock='1';
  address<=X"0000005B";
  write_data<= X"00000143";
  wait until clock'event and clock='1';
  address<=X"0000005C";
  write_data<=X"00000144";
  wait until clock'event and clock='1';
  address<=X"0000005D";
  write_data<= X"00000145";
  wait until clock'event and clock='1';
  address<=X"0000005E";
  write_data<= X"00000146";
  wait until clock'event and clock='1';
  address<=X"0000005F";
  write_data<=X"00000147";
  wait until clock'event and clock='1';
  address<=X"00000060";
  write_data<= X"00000148";
  wait until clock'event and clock='1';
  address<=X"00000061";
  write_data<= X"00000149";
  wait until clock'event and clock='1';
  address<=X"00000062";
  write_data<=X"00000150";
  wait until clock'event and clock='1';
  address<=X"00000063";
  write_data<= X"00000151";
  wait until clock'event and clock='1';
  address<=X"00000064";
  write_data<= X"00000152";
  wait until clock'event and clock='1';
  address<=X"00000065";
  write_data<= X"00000153";
  wait until clock'event and clock='1';
  address<=X"00000066";
  write_data<=X"00000154";
  wait until clock'event and clock='1';
  address<=X"00000067";
  write_data<= X"00000155";
  wait until clock'event and clock='1';
  address<=X"00000068";
  write_data<= X"00000156";
  wait until clock'event and clock='1';
  address<=X"00000069";
  write_data<=X"00000157";
  wait until clock'event and clock='1';
  address<=X"0000006A";
  write_data<= X"00000158";
  wait until clock'event and clock='1';
  address<=X"0000006B";
  write_data<= X"00000159";
  wait until clock'event and clock='1';
  address<=X"0000006C";
  write_data<=X"00000160";
  wait until clock'event and clock='1';
  address<=X"0000006D";
  write_data<= X"00000161";
  wait until clock'event and clock='1';
  address<=X"0000006E";
  write_data<= X"00000162";
  wait until clock'event and clock='1';
  address<=X"0000006F";
  write_data<= X"00000163";
  wait until clock'event and clock='1';
  address<=X"00000070";
  write_data<=X"00000164";
  wait until clock'event and clock='1';
  address<=X"00000071";
  write_data<= X"00000165";
  wait until clock'event and clock='1';
  address<=X"00000072";
  write_data<= X"00000166";
  wait until clock'event and clock='1';
  address<=X"00000073";
  write_data<=X"00000167";
  wait until clock'event and clock='1';
  address<=X"00000074";
  write_data<= X"00000168";
  wait until clock'event and clock='1';
  address<=X"00000075";
  write_data<= X"00000169";
  wait until clock'event and clock='1';
  address<=X"00000076";
  write_data<=X"00000170";
  wait until clock'event and clock='1';
  address<=X"00000077";
  write_data<= X"00000171";
  wait until clock'event and clock='1';
  address<=X"00000078";
  write_data<= X"00000172";
  wait until clock'event and clock='1';
  address<=X"00000079";
  write_data<= X"00000173";
  wait until clock'event and clock='1';
  address<=X"0000007A";
  write_data<=X"00000174";
  wait until clock'event and clock='1';
  address<=X"0000007B";
  write_data<= X"00000175";
  wait until clock'event and clock='1';
  address<=X"0000007C";
  write_data<= X"00000176";
  wait until clock'event and clock='1';
  address<=X"0000007D";
  write_data<=X"00000177";
  wait until clock'event and clock='1';
  address<=X"0000007E";
  write_data<= X"00000178";
  wait until clock'event and clock='1';
  address<=X"0000007F";
  write_data<= X"00000179";
  wait until clock'event and clock='1';
  address<=X"00000080";
  write_data<=X"00000180";
  wait until clock'event and clock='1';
  address<=X"00000081";
  write_data<= X"00000181";
  wait until clock'event and clock='1';
  address<=X"00000082";
  write_data<= X"00000182";
  wait until clock'event and clock='1';
  address<=X"00000083";
  write_data<= X"00000183";
  wait until clock'event and clock='1';
  address<=X"00000084";
  write_data<=X"00000184";
  wait until clock'event and clock='1';
  address<=X"00000085";
  write_data<= X"00000185";
  wait until clock'event and clock='1';
  address<=X"00000086";
  write_data<= X"00000186";
  wait until clock'event and clock='1';
  address<=X"00000087";
  write_data<=X"00000187";
  wait until clock'event and clock='1';
  address<=X"00000088";
  write_data<= X"00000188";
  wait until clock'event and clock='1';
  address<=X"00000089";
  write_data<= X"00000189";
  wait until clock'event and clock='1';
  address<=X"0000008A";
write_data<=X"00000190" ;
wait until clock'event and clock='1';
  address<=X"0000008B";
write_data<=X"00000191";
wait until clock'event and clock='1';
  address<=X"0000008C";
write_data<= X"00000192";
wait until clock'event and clock='1';
  address<=X"0000008D";
write_data<= X"00000193";
wait until clock'event and clock='1';
  address<=X"0000008E";
write_data<=X"00000194";
wait until clock'event and clock='1';
  address<=X"0000008F";
write_data<= X"00000195";
wait until clock'event and clock='1';
  address<=X"00000090";
write_data<= X"00000196";
wait until clock'event and clock='1';
  address<=X"00000091";
write_data<=X"00000197";
wait until clock'event and clock='1';
  address<=X"00000092";
write_data<= X"00000198";
---------
wait until clock'event and clock='1';
  address<=X"00000093";
write_data<= X"00000199";
wait until clock'event and clock='1';
  address<=X"00000094";
write_data<=X"00000200";
wait until clock'event and clock='1';
  address<=X"00000095";
write_data<= X"00000201";
wait until clock'event and clock='1';
  address<=X"00000096";
write_data<= X"00000202";
wait until clock'event and clock='1';
  address<=X"00000097";
write_data<= X"00000203";
wait until clock'event and clock='1';
  address<=X"00000098";
write_data<=X"00000204";
wait until clock'event and clock='1';
  address<=X"00000099";
write_data<= X"00000205";
wait until clock'event and clock='1';
  address<=X"0000009A";
write_data<= X"00000206";
wait until clock'event and clock='1';
  address<=X"0000009B";
write_data<=X"00000207";
wait until clock'event and clock='1';
  address<=X"0000009C";
write_data<=X"00000208";
wait until clock'event and clock='1';
  address<=X"0000009D";
write_data<=X"00000209";
wait until clock'event and clock='1';
  address<=X"0000009E";
write_data<=X"00000210";
wait until clock'event and clock='1';
  address<=X"0000009F";
write_data<= X"00000211";
wait until clock'event and clock='1';
  address<=X"000000A0";
write_data<= X"00000212";
wait until clock'event and clock='1';
  address<=X"000000A1";
write_data<= X"00000213";
wait until clock'event and clock='1';
  address<=X"000000A2";
write_data<=X"00000214";
wait until clock'event and clock='1';
  address<=X"000000A3";
write_data<=X"00000215";
wait until clock'event and clock='1';
  address<=X"000000A4";
write_data<= X"00000216";
wait until clock'event and clock='1';
  address<=X"000000A5";
write_data<=X"00000217";
wait until clock'event and clock='1';
  address<=X"000000A6";
write_data<=X"00000218";
wait until clock'event and clock='1';
  address<=X"000000A7";
write_data<= X"00000219";
wait until clock'event and clock='1';
  address<=X"000000A8";
write_data<=X"00000220";
wait until clock'event and clock='1';
  address<=X"000000A9";
write_data<= X"00000221";
wait until clock'event and clock='1';
  address<=X"000000AA";
write_data<= X"00000222";
wait until clock'event and clock='1';
  address<=X"000000AB";
write_data<= X"00000223";
wait until clock'event and clock='1';
  address<=X"000000AC";
write_data<=X"00000224";
wait until clock'event and clock='1';
  address<=X"000000AD";
write_data<=X"00000225";
wait until clock'event and clock='1';
  address<=X"000000AE";
write_data<=X"00000226";
wait until clock'event and clock='1';
  address<=X"000000AF";
write_data<=X"00000227";
wait until clock'event and clock='1';
  address<=X"000000B0";
write_data<= X"00000228";
wait until clock'event and clock='1';
  address<=X"000000B1";
write_data<= X"00000229";
wait until clock'event and clock='1';
  address<=X"000000B2";
write_data<=X"00000230";
wait until clock'event and clock='1';
  address<=X"000000B3";
write_data<=X"00000231";
wait until clock'event and clock='1';
  address<=X"000000B4";
write_data<=X"00000232";
wait until clock'event and clock='1';
  address<=X"000000B5";
write_data<=X"00000233";
wait until clock'event and clock='1';
  address<=X"000000B6";
write_data<=X"00000234";
wait until clock'event and clock='1';
  address<=X"000000B7";
write_data<= X"00000235";
wait until clock'event and clock='1';
  address<=X"000000B8";
write_data<= X"00000236";
wait until clock'event and clock='1';
  address<=X"000000B9";
write_data<=X"00000237";
wait until clock'event and clock='1';
  address<=X"000000BA";
write_data<=X"00000238";
wait until clock'event and clock='1';
  address<=X"000000BB";
write_data<=X"00000239";
wait until clock'event and clock='1';
  address<=X"000000BC";
write_data<=X"00000240";
wait until clock'event and clock='1';
  address<=X"000000BD";
write_data<= X"00000241";
wait until clock'event and clock='1';
  address<=X"000000BE";
write_data<= X"00000242";
wait until clock'event and clock='1';
  address<=X"000000BF";
write_data<= X"00000243";
wait until clock'event and clock='1';
  address<=X"000000C0";
write_data<= X"00000244";
wait until clock'event and clock='1';
  address<=X"000000C1";
write_data<= X"00000245";
wait until clock'event and clock='1';
  address<=X"000000C2";
write_data<= X"00000246";
wait until clock'event and clock='1';
  address<=X"000000C3";
write_data<=X"00000247";
wait until clock'event and clock='1';
  address<=X"000000C4";
write_data<=X"00000248";
wait until clock'event and clock='1';
  address<=X"000000C5";
write_data<=X"00000249";
wait until clock'event and clock='1';
  address<=X"000000C6";
write_data<=X"00000250";
wait until clock'event and clock='1';
  address<=X"000000C7";
write_data<= X"00000251";
wait until clock'event and clock='1';
  address<=X"000000C8";
write_data<= X"00000252";
wait until clock'event and clock='1';
  address<=X"000000C9";
write_data<= X"00000253";
wait until clock'event and clock='1';
  address<=X"000000CA";
write_data<=X"00000254";
wait until clock'event and clock='1';
  address<=X"000000CB";
write_data<=X"00000255";
wait until clock'event and clock='1';
  address<=X"000000CC";
write_data<= X"00000256";
wait until clock'event and clock='1';
  address<=X"000000CD";
write_data<=X"00000257";
wait until clock'event and clock='1';
  address<=X"000000CE";
write_data<=X"00000258";
wait until clock'event and clock='1';
  address<=X"000000CF";
write_data<=X"00000259";
wait until clock'event and clock='1';
  address<=X"000000D0";
write_data<=X"00000260";
wait until clock'event and clock='1';
  address<=X"000000D1";
write_data<= X"00000261";
wait until clock'event and clock='1';
  address<=X"000000D2";
write_data<= X"00000262";
wait until clock'event and clock='1';
  address<=X"000000D3";
write_data<=X"00000263";
wait until clock'event and clock='1';
  address<=X"000000D4";
write_data<=X"00000264";
wait until clock'event and clock='1';
  address<=X"000000D5";
write_data<= X"00000265";
wait until clock'event and clock='1';
  address<=X"000000D6";
write_data<= X"00000266";
wait until clock'event and clock='1';
  address<=X"000000D7";
write_data<=X"00000267";
wait until clock'event and clock='1';
  address<=X"000000D8";
write_data<=X"00000268";
wait until clock'event and clock='1';
  address<=X"000000D9";
write_data<=X"00000269";
wait until clock'event and clock='1';
  address<=X"000000DA";
write_data<=X"00000270";
wait until clock'event and clock='1';
  address<=X"000000DB";
write_data<= X"00000271";
wait until clock'event and clock='1';
  address<=X"000000DC";
write_data<= X"00000272";
wait until clock'event and clock='1';
  address<=X"000000DD";
write_data<= X"00000273";
wait until clock'event and clock='1';
  address<=X"000000DE";
write_data<=X"00000274";
wait until clock'event and clock='1';
  address<=X"000000DF";
write_data<=X"00000275";
wait until clock'event and clock='1';
  address<=X"000000E0";
write_data<=X"00000276";
wait until clock'event and clock='1';
  address<=X"000000E1";
write_data<=X"00000277";
wait until clock'event and clock='1';
  address<=X"000000E2";
write_data<=X"00000278";
wait until clock'event and clock='1';
  address<=X"000000E3";
write_data<= X"00000279";
wait until clock'event and clock='1';
  address<=X"000000E4";
write_data<=X"00000280";
wait until clock'event and clock='1';
  address<=X"000000E5";
write_data<= X"00000281";
wait until clock'event and clock='1';
  address<=X"000000E6";
write_data<=X"00000282";
wait until clock'event and clock='1';
  address<=X"000000E7";
write_data<= X"00000283";
wait until clock'event and clock='1';
  address<=X"000000E8";
write_data<=X"00000284";
wait until clock'event and clock='1';
  address<=X"000000E9";
write_data<=X"00000285";
wait until clock'event and clock='1';
  address<=X"000000EA";
write_data<=X"00000286";
wait until clock'event and clock='1';
  address<=X"000000EB";
write_data<=X"00000287";
wait until clock'event and clock='1';
  address<=X"000000EC";
write_data<= X"00000288";
wait until clock'event and clock='1';
  address<=X"000000ED";
write_data<= X"00000289";
wait until clock'event and clock='1';
  address<=X"000000EE";
write_data<=X"00000290";
wait until clock'event and clock='1';
  address<=X"000000EF";
write_data<= X"00000291";
wait until clock'event and clock='1';
  address<=X"000000F0";
write_data<= X"00000292";
wait until clock'event and clock='1';
  address<=X"000000F1";
write_data<=X"00000293";
wait until clock'event and clock='1';
  address<=X"000000F2";
write_data<=X"00000294";
wait until clock'event and clock='1';
  address<=X"000000F3";
write_data<= X"00000295";
wait until clock'event and clock='1';
  address<=X"000000F4";
write_data<= X"00000296";
wait until clock'event and clock='1';
  address<=X"000000F5";
write_data<=X"00000297";
wait until clock'event and clock='1';
  address<=X"000000F6";
write_data<=X"00000298";
wait until clock'event and clock='1';
  address<=X"000000F7";
write_data<=X"00000299";
wait until clock'event and clock='1';
  address<=X"000000F8";
write_data<=X"00000300";
wait until clock'event and clock='1';
  address<=X"000000F9";
write_data<=X"00000301";
wait until clock'event and clock='1';
  address<=X"000000FA";
write_data<=X"00000302";
wait until clock'event and clock='1';
  address<=X"000000FB";
write_data<= X"00000303";
wait until clock'event and clock='1';
  address<=X"000000FC";
write_data<=X"00000304";
wait until clock'event and clock='1';
  address<=X"000000FD";
write_data<=X"00000305";
wait until clock'event and clock='1';
  address<=X"000000FE";
write_data<=X"00000306";
wait until clock'event and clock='1';
  address<=X"000000FF";
write_data<=X"00000307";
wait until clock'event and clock='1';
  address<=X"00000100";
write_data<= X"00000308";
wait until clock'event and clock='1';
  address<=X"00000101";
write_data<= X"00000309";
wait until clock'event and clock='1';
  address<=X"00000102";
write_data<=X"00000310";
wait until clock'event and clock='1';
  address<=X"00000103";
write_data<= X"00000311";
wait until clock'event and clock='1';
  address<=X"00000104";
write_data<= X"00000312";
wait until clock'event and clock='1';
  address<=X"00000105";
write_data<= X"00000313";
wait until clock'event and clock='1';
  address<=X"00000106";
write_data<=X"00000314";
wait until clock'event and clock='1';
  address<=X"00000107";
write_data<= X"00000315";
wait until clock'event and clock='1';
  address<=X"00000108";
write_data<= X"00000316";
wait until clock'event and clock='1';
  address<=X"00000109";
write_data<=X"00000317";
wait until clock'event and clock='1';
  address<=X"0000010A";
write_data<=X"00000318";
wait until clock'event and clock='1';
  address<=X"0000010B";
write_data<=X"00000319";
wait until clock'event and clock='1';
  address<=X"0000010C";
write_data<=X"00000320";
wait until clock'event and clock='1';
  address<=X"0000010D";
write_data<= X"00000321";
wait until clock'event and clock='1';
  address<=X"0000010E";
write_data<= X"00000322";
wait until clock'event and clock='1';
  address<=X"0000010F";
write_data<= X"00000323";
wait until clock'event and clock='1';
  address<=X"00000110";
write_data<=X"00000324";
wait until clock'event and clock='1';
  address<=X"00000111";
write_data<= X"00000325";
wait until clock'event and clock='1';
  address<=X"00000112";
write_data<= X"00000326";
wait until clock'event and clock='1';
  address<=X"00000113";
write_data<=X"00000327";
wait until clock'event and clock='1';
  address<=X"00000114";
write_data<=X"00000328";
wait until clock'event and clock='1';
  address<=X"00000115";
write_data<= X"00000329";
wait until clock'event and clock='1';
  address<=X"00000116";
write_data<=X"00000330";
wait until clock'event and clock='1';
  address<=X"00000117";
write_data<= X"00000331";
wait until clock'event and clock='1';
  address<=X"00000118";
write_data<= X"00000332";
wait until clock'event and clock='1';
  address<=X"00000119";
write_data<= X"00000333";
wait until clock'event and clock='1';
  address<=X"0000011A";
write_data<=X"00000334";
wait until clock'event and clock='1';
  address<=X"0000011B";
write_data<=X"00000335";
wait until clock'event and clock='1';
  address<=X"0000011C";
write_data<=X"00000336";
wait until clock'event and clock='1';
  address<=X"0000011D";
write_data<=X"00000337";
wait until clock'event and clock='1';
  address<=X"0000011E";
write_data<= X"00000338";
wait until clock'event and clock='1';
  address<=X"0000011F";
write_data<= X"00000339";
wait until clock'event and clock='1';
  address<=X"00000120";
write_data<=X"00000340";
wait until clock'event and clock='1';
  address<=X"00000121";
write_data<= X"00000341";
wait until clock'event and clock='1';
  address<=X"00000122";
write_data<= X"00000342";
wait until clock'event and clock='1';
  address<=X"00000123";
write_data<= X"00000343";
wait until clock'event and clock='1';
  address<=X"00000124";
write_data<=X"00000344";
wait until clock'event and clock='1';
  address<=X"00000125";
write_data<=X"00000345";
wait until clock'event and clock='1';
  address<=X"00000126";
write_data<=X"00000346";
wait until clock'event and clock='1';
  address<=X"00000127";
write_data<=X"00000347";
wait until clock'event and clock='1';
  address<=X"00000128";
write_data<= X"00000348";
wait until clock'event and clock='1';
  address<=X"00000129";
write_data<= X"00000349";
wait until clock'event and clock='1';
  address<=X"0000012A";
write_data<=X"00000350";
wait until clock'event and clock='1';
  address<=X"0000012B";
write_data<= X"00000351";
wait until clock'event and clock='1';
  address<=X"0000012C";
write_data<= X"00000352";
wait until clock'event and clock='1';
  address<=X"0000012D";
write_data<= X"00000353";
wait until clock'event and clock='1';
  address<=X"0000012E";
write_data<=X"00000354";
wait until clock'event and clock='1';
  address<=X"0000012F";
write_data<=X"00000355";
wait until clock'event and clock='1';
  address<=X"00000130";
write_data<=X"00000356";
wait until clock'event and clock='1';
  address<=X"00000131";
write_data<=X"00000357";
wait until clock'event and clock='1';
  address<=X"00000132";
write_data<= X"00000358";
wait until clock'event and clock='1';
  address<=X"00000133";
write_data<= X"00000359";
wait until clock'event and clock='1';
  address<=X"00000134";
write_data<=X"00000360";
wait until clock'event and clock='1';
  address<=X"00000135";
write_data<= X"00000361";
wait until clock'event and clock='1';
  address<=X"00000136";
write_data<= X"00000362";
wait until clock'event and clock='1';
  address<=X"00000137";
write_data<= X"00000363";
wait until clock'event and clock='1';
  address<=X"00000138";
write_data<=X"00000364";
wait until clock'event and clock='1';
  address<=X"00000139";
write_data<= X"00000365";
wait until clock'event and clock='1';
  address<=X"0000013A";
write_data<= X"00000366";
wait until clock'event and clock='1';
  address<=X"0000013B";
write_data<=X"00000367";
wait until clock'event and clock='1';
  address<=X"0000013C";
write_data<=X"00000368";
wait until clock'event and clock='1';
  address<=X"0000013D";
write_data<=X"00000369";
wait until clock'event and clock='1';
  address<=X"0000013E";
write_data<=X"00000370";
wait until clock'event and clock='1';
  address<=X"0000013F";
write_data<=X"00000371";
wait until clock'event and clock='1';
  address<=X"00000140";
write_data<=X"00000372";
wait until clock'event and clock='1';
  address<=X"00000141";
write_data<=X"00000373";
wait until clock'event and clock='1';
  address<=X"00000142";
write_data<=X"00000374";
wait until clock'event and clock='1';
  address<=X"00000143";
write_data<= X"00000375";
wait until clock'event and clock='1';
  address<=X"00000144";
write_data<= X"00000376";
wait until clock'event and clock='1';
  address<=X"00000145";
write_data<=X"00000377";
wait until clock'event and clock='1';
  address<=X"00000146";
write_data<= X"00000378";
wait until clock'event and clock='1';
  address<=X"00000147";
write_data<= X"00000379";
wait until clock'event and clock='1';
  address<=X"00000148";
write_data<=X"00000380";
wait until clock'event and clock='1';
  address<=X"00000149";
write_data<= X"00000381";
wait until clock'event and clock='1';
  address<=X"0000014A";
write_data<= X"00000382";
wait until clock'event and clock='1';
  address<=X"0000014B";
write_data<=X"00000383";
wait until clock'event and clock='1';
  address<=X"0000014C";
write_data<=X"00000384";
wait until clock'event and clock='1';
  address<=X"0000014D";
write_data<= X"00000385";
wait until clock'event and clock='1';
  address<=X"0000014E";
write_data<= X"00000386";
wait until clock'event and clock='1';
  address<=X"0000014F";
write_data<=X"00000387";
wait until clock'event and clock='1';
  address<=X"00000150";
write_data<=X"00000388";
wait until clock'event and clock='1';
  address<=X"00000151";
write_data<=X"00000389";
wait until clock'event and clock='1';
  address<=X"00000152";
write_data<=X"00000390";
wait until clock'event and clock='1';
  address<=X"00000153";
write_data<= X"00000391";
wait until clock'event and clock='1';
  address<=X"00000154";
write_data<= X"00000392";
wait until clock'event and clock='1';
  address<=X"00000155";
write_data<= X"00000393";
wait until clock'event and clock='1';
  address<=X"00000156";
write_data<=X"00000394";
wait until clock'event and clock='1';
  address<=X"00000157";
write_data<=X"00000395";
wait until clock'event and clock='1';
  address<=X"00000158";
write_data<=X"00000396";
wait until clock'event and clock='1';
  address<=X"00000159";
write_data<=X"00000397";
wait until clock'event and clock='1';
  address<=X"0000015A";
write_data<= X"00000398";
wait until clock'event and clock='1';
  address<=X"0000015B";
write_data<= X"00000399";
wait until clock'event and clock='1';
  address<=X"0000015C";
write_data<=X"00000400";
wait until clock'event and clock='1';
  address<=X"0000015D";
write_data<=X"00000401";
wait until clock'event and clock='1';
  address<=X"0000015E";
write_data<= X"00000402";
wait until clock'event and clock='1';
  address<=X"0000015F";
write_data<= X"00000403";
wait until clock'event and clock='1';
  address<=X"00000160";
write_data<=X"00000404";
wait until clock'event and clock='1';
  address<=X"00000161";
write_data<=X"00000405";
wait until clock'event and clock='1';
  address<=X"00000162";
write_data<=X"00000406";
wait until clock'event and clock='1';
  address<=X"00000163";
write_data<=X"00000407";
wait until clock'event and clock='1';
  address<=X"00000164";
write_data<= X"00000408";
wait until clock'event and clock='1';
  address<=X"00000165";
write_data<=X"00000409";
wait until clock'event and clock='1';
  address<=X"00000166";
write_data<=X"00000410";
wait until clock'event and clock='1';
  address<=X"00000167";
write_data<= X"00000411";
wait until clock'event and clock='1';
  address<=X"00000168";
write_data<= X"00000412";
wait until clock'event and clock='1';
  address<=X"00000169";
write_data<= X"00000413";
wait until clock'event and clock='1';
  address<=X"0000016A";
write_data<=X"00000414";
wait until clock'event and clock='1';
  address<=X"0000016B";
write_data<= X"00000415";
wait until clock'event and clock='1';
  address<=X"0000016C";
write_data<= X"00000416";
wait until clock'event and clock='1';
  address<=X"0000016D";
write_data<=X"00000417";
wait until clock'event and clock='1';
  address<=X"0000016E";
write_data<= X"00000418";
wait until clock'event and clock='1';
  address<=X"0000016F";
write_data<= X"00000419";
wait until clock'event and clock='1';
  address<=X"00000170";
write_data<=X"00000420";
wait until clock'event and clock='1';
  address<=X"00000171";
write_data<=X"00000421";
wait until clock'event and clock='1';
  address<=X"00000172";
write_data<= X"00000422";
wait until clock'event and clock='1';
  address<=X"00000173";
write_data<= X"00000423";
wait until clock'event and clock='1';
  address<=X"00000174";
write_data<=X"00000424";
wait until clock'event and clock='1';
  address<=X"00000175";
write_data<= X"00000425";
wait until clock'event and clock='1';
  address<=X"00000176";
write_data<= X"00000426";
wait until clock'event and clock='1';
  address<=X"00000177";
write_data<=X"00000427";
wait until clock'event and clock='1';
  address<=X"00000178";
write_data<= X"00000428";
wait until clock'event and clock='1';
  address<=X"00000179";
write_data<=X"00000429";
wait until clock'event and clock='1';
  address<=X"0000017A";
write_data<=X"00000430";
wait until clock'event and clock='1';
  address<=X"0000017B";
write_data<= X"00000431";
wait until clock'event and clock='1';
  address<=X"0000017C";
write_data<= X"00000432";
wait until clock'event and clock='1';
  address<=X"0000017D";
write_data<= X"00000433";
wait until clock'event and clock='1';
  address<=X"0000017E";
write_data<=X"00000434";
wait until clock'event and clock='1';
  address<=X"0000017F";
write_data<= X"00000435";
wait until clock'event and clock='1';
  address<=X"00000180";
write_data<= X"00000436";
wait until clock'event and clock='1';
  address<=X"00000181";
write_data<=X"00000437";
wait until clock'event and clock='1';
  address<=X"00000182";
write_data<= X"00000438" ;
wait until clock'event and clock='1';
  address<=X"00000183";
write_data<=X"00000439";
wait until clock'event and clock='1';
  address<=X"00000184";
write_data<=X"00000440";
wait until clock'event and clock='1';
  address<=X"00000185";
write_data<= X"00000441";
wait until clock'event and clock='1';
  address<=X"00000186";
write_data<= X"00000442";
wait until clock'event and clock='1';
  address<=X"00000187";
write_data<= X"00000443";
wait until clock'event and clock='1';
  address<=X"00000188";
write_data<=X"00000444";
wait until clock'event and clock='1';
  address<=X"00000189";
write_data<= X"00000445";
wait until clock'event and clock='1';
  address<=X"0000018A";
write_data<= X"00000446";
wait until clock'event and clock='1';
  address<=X"0000018B";
write_data<=X"00000447";
wait until clock'event and clock='1';
  address<=X"0000018C";
write_data<= X"00000448";
wait until clock'event and clock='1';
  address<=X"0000018D";
write_data<= X"00000449";
wait until clock'event and clock='1';
  address<=X"0000018E";
write_data<=X"00000450";
wait until clock'event and clock='1';
  address<=X"0000018F";
write_data<= X"00000451";
wait until clock'event and clock='1';
  address<=X"00000190";
write_data<= X"00000452";
wait until clock'event and clock='1';
  address<=X"00000191";
write_data<= X"00000453";
wait until clock'event and clock='1';
  address<=X"00000192";
write_data<=X"00000454";
wait until clock'event and clock='1';
  address<=X"00000193";
write_data<= X"00000455";
wait until clock'event and clock='1';
  address<=X"00000194";
write_data<= X"00000456";
wait until clock'event and clock='1';
  address<=X"00000195";
write_data<=X"00000457";
wait until clock'event and clock='1';
  address<=X"00000196";
write_data<= X"00000458";
wait until clock'event and clock='1';
  address<=X"00000197";
write_data<= X"00000459";
wait until clock'event and clock='1';
  address<=X"00000198";
write_data<=X"00000460";
wait until clock'event and clock='1';
  address<=X"00000199";
write_data<= X"00000461";
wait until clock'event and clock='1';
  address<=X"0000019A";
write_data<= X"00000462";
wait until clock'event and clock='1';
  address<=X"0000019B";
write_data<= X"00000463";
wait until clock'event and clock='1';
  address<=X"0000019C";
write_data<=X"00000464";
wait until clock'event and clock='1';
  address<=X"0000019D";
write_data<= X"00000465";
wait until clock'event and clock='1';
  address<=X"0000010E";
write_data<= X"00000466";
wait until clock'event and clock='1';
  address<=X"0000019F";
write_data<=X"00000467";
wait until clock'event and clock='1';
  address<=X"000001A0";
write_data<= X"00000468";
wait until clock'event and clock='1';
  address<=X"000001A1";
write_data<= X"00000469";
wait until clock'event and clock='1';
  address<=X"000001A2";
write_data<=X"00000470";
wait until clock'event and clock='1';
  address<=X"000001A3";
write_data<= X"00000471";
wait until clock'event and clock='1';
  address<=X"00000143";
write_data<= X"00000472";
wait until clock'event and clock='1';
  address<=X"000001A5";
write_data<= X"00000473";
wait until clock'event and clock='1';
  address<=X"000001A6";
write_data<=X"00000474";
wait until clock'event and clock='1';
  address<=X"000001A7";
write_data<= X"00000475";
wait until clock'event and clock='1';
  address<=X"000001A8";
write_data<= X"00000476";
wait until clock'event and clock='1';
  address<=X"000001A9";
write_data<=X"00000477";
wait until clock'event and clock='1';
  address<=X"000001AA";
write_data<= X"00000478";
wait until clock'event and clock='1';
  address<=X"000001AB";
write_data<= X"00000479";
wait until clock'event and clock='1';
  address<=X"000001AC";
write_data<=X"00000480";
wait until clock'event and clock='1';
  address<=X"000001AD";
write_data<= X"00000481";
wait until clock'event and clock='1';
  address<=X"000001AE";
write_data<= X"00000482";
wait until clock'event and clock='1';
  address<=X"000001AF";
write_data<= X"00000483";
wait until clock'event and clock='1';
  address<=X"000001B0";
write_data<=X"00000484";
wait until clock'event and clock='1';
  address<=X"000001B1";
write_data<= X"00000485";
wait until clock'event and clock='1';
  address<=X"000001B2";
write_data<= X"00000486";
wait until clock'event and clock='1';
  address<=X"000001B3";
write_data<=X"00000487";
wait until clock'event and clock='1';
  address<=X"000001B4";
write_data<= X"00000488";
wait until clock'event and clock='1';
  address<=X"000001B5";
write_data<= X"00000489";
wait until clock'event and clock='1';
  address<=X"000001B6";
write_data<=X"00000490";
wait until clock'event and clock='1';
  address<=X"000001B7";
write_data<= X"00000491";
wait until clock'event and clock='1';
  address<=X"000001B8";
write_data<= X"00000492";
wait until clock'event and clock='1';
  address<=X"000001B9";
write_data<= X"00000493";
wait until clock'event and clock='1';
  address<=X"000001BA";
write_data<=X"00000494";
wait until clock'event and clock='1';
  address<=X"000001BB";
write_data<= X"00000495";
wait until clock'event and clock='1';
  address<=X"000001BC";
write_data<= X"00000496";
wait until clock'event and clock='1';
  address<=X"000001BD";
write_data<=X"00000497";
wait until clock'event and clock='1';
  address<=X"000001BE";
write_data<= X"00000498";
wait until clock'event and clock='1';
  address<=X"000001BF";
write_data<= X"00000499";
wait until clock'event and clock='1';
  address<=X"000001C0";
write_data<=X"00000500";
wait until clock'event and clock='1';
  address<=X"000001C1";
write_data<= X"00000501";
wait until clock'event and clock='1';
  address<=X"000001C2";
write_data<= X"00000502";
wait until clock'event and clock='1';
  address<=X"000001C3";
write_data<= X"00000503";
wait until clock'event and clock='1';
  address<=X"000001C4";
write_data<=X"00000504";
wait until clock'event and clock='1';
  address<=X"000001C5";
write_data<= X"00000505";
wait until clock'event and clock='1';
  address<=X"000001C6";
write_data<= X"00000506";
wait until clock'event and clock='1';
  address<=X"000001C7";
write_data<=X"00000507";
wait until clock'event and clock='1';
  address<=X"000001C8";
write_data<= X"00000508";
wait until clock'event and clock='1';
  address<=X"000001C9";
write_data<= X"00000509";
wait until clock'event and clock='1';
  address<=X"000001CA";
write_data<=X"00000510";
wait until clock'event and clock='1';
  address<=X"000001CB";
write_data<= X"00000511";
wait until clock'event and clock='1';
  address<=X"000001CC";
write_data<= X"00000512";
wait until clock'event and clock='1';
  address<=X"000001CD";
write_data<= X"00000513";
wait until clock'event and clock='1';
  address<=X"000001CE";
write_data<=X"00000514";
wait until clock'event and clock='1';
  address<=X"000001CF";
write_data<= X"00000515";
wait until clock'event and clock='1';
  address<=X"000001D0";
write_data<= X"00000516";
wait until clock'event and clock='1';
  address<=X"000001D1";
write_data<=X"00000517";
wait until clock'event and clock='1';
  address<=X"000001D2";
write_data<= X"00000518";
wait until clock'event and clock='1';
  address<=X"000001D3";
write_data<= X"00000519";
wait until clock'event and clock='1';
  address<=X"000001D4";
write_data<=X"00000520";
wait until clock'event and clock='1';
  address<=X"000001D5";
write_data<= X"00000521";
wait until clock'event and clock='1';
  address<=X"000001D6";
write_data<= X"00000522";
wait until clock'event and clock='1';
  address<=X"000001D7";
write_data<= X"00000523";
wait until clock'event and clock='1';
  address<=X"000001D8";
write_data<=X"00000524";
wait until clock'event and clock='1';
  address<=X"000001D9";
write_data<= X"00000525";
wait until clock'event and clock='1';
  address<=X"000001DA";
write_data<= X"00000526";
wait until clock'event and clock='1';
  address<=X"000001DB";
write_data<=X"00000527";
wait until clock'event and clock='1';
  address<=X"000001DC";
write_data<= X"00000528";
wait until clock'event and clock='1';
  address<=X"000001DD";
write_data<= X"00000529";
wait until clock'event and clock='1';
  address<=X"000001DE";
write_data<=X"00000530";
wait until clock'event and clock='1';
  address<=X"000001DF";
write_data<= X"00000531";
wait until clock'event and clock='1';
  address<=X"000001E0";
write_data<= X"00000532";
wait until clock'event and clock='1';
  address<=X"000001E1";
write_data<= X"00000533";
wait until clock'event and clock='1';
  address<=X"000001E2";
write_data<=X"00000534";
wait until clock'event and clock='1';
  address<=X"000001E3";
write_data<= X"00000535";
wait until clock'event and clock='1';
  address<=X"000001E4";
write_data<= X"00000536";
wait until clock'event and clock='1';
  address<=X"000001E5";
write_data<=X"00000537";
wait until clock'event and clock='1';
  address<=X"000001E6";
write_data<= X"00000538";
wait until clock'event and clock='1';
  address<=X"000001E7";
write_data<= X"00000539";
wait until clock'event and clock='1';
  address<=X"000001E8";
write_data<=X"00000540";
wait until clock'event and clock='1';
  address<=X"000001E9";
write_data<= X"00000541";
wait until clock'event and clock='1';
  address<=X"000001EA";
write_data<= X"00000542";
wait until clock'event and clock='1';
  address<=X"000001EB";
write_data<= X"00000543";
wait until clock'event and clock='1';
  address<=X"000001EC";
write_data<=X"00000544";
wait until clock'event and clock='1';
  address<=X"000001ED";
write_data<= X"00000545";
wait until clock'event and clock='1';
  address<=X"000001EE";
write_data<= X"00000546";
wait until clock'event and clock='1';
  address<=X"000001EF";
write_data<=X"00000547";
wait until clock'event and clock='1';
  address<=X"000001F0";
write_data<= X"00000548";
wait until clock'event and clock='1';
  address<=X"000001F1";
write_data<= X"00000549";
wait until clock'event and clock='1';
  address<=X"000001F2";
write_data<=X"00000550";
wait until clock'event and clock='1';
  address<=X"000001F3";
write_data<= X"00000551";
wait until clock'event and clock='1';
  address<=X"000001F4";
write_data<=X"00000552";
wait until clock'event and clock='1';
  address<=X"000001F5";
write_data<= X"00000553";
wait until clock'event and clock='1';
  address<=X"000001F6";
write_data<=X"00000554";
wait until clock'event and clock='1';
  address<=X"000001F7";
write_data<= X"00000555";
wait until clock'event and clock='1';
  address<=X"000001F8";
write_data<= X"00000556";
wait until clock'event and clock='1';
  address<=X"000001F9";
write_data<=X"00000557";
wait until clock'event and clock='1';
  address<=X"000001FA";
write_data<= X"00000558";
wait until clock'event and clock='1';
  address<=X"000001FB";
write_data<= X"00000559";
wait until clock'event and clock='1';
  address<=X"000001FC";
write_data<=X"00000560";
wait until clock'event and clock='1';
  address<=X"000001FD";
write_data<= X"00000561";
wait until clock'event and clock='1';
  address<=X"000001FE";
write_data<= X"00000562"; 
wait until clock'event and clock='1';
  address<=X"000001FF";
write_data<=X"00000563"; 
wait until clock'event and clock='1';
  end process;
end;
